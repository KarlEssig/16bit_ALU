module ShiftRight(input [15:0] a, b, output [15:0] s);
	assign res = a >> b;
endmodule
